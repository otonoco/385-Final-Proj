module mario_s (
        input Reset, frame_clk, Clk,
        input [31:0] keycode,
        input [9:0] DrawX, DrawY,
        input mario_alive,

        input [23:0] mario_sl, mario_sr, mario_rl1, mario_rl2, mario_rl3, mario_rr1, mario_rr2, mario_rr3, mario_jr, mario_jl, mario_die,

        output logic [9:0] mario_x, mario_y, process, mario_y_motion,
        output logic mario, mario_in_air,
        output logic [23:0] mario_counter, 
        output logic [23:0] mario_pic_out
);
    logic w, s, a, d;
    logic sl, sr, rr1, rr2, rr3, rl1, rl2, rl3, jr, jl, il, ir, gr, gl, di;

    assign a = ((keycode[15:8] == 8'h04) | (keycode[7:0] == 8'h04)|(keycode[23:16] == 8'h04) | (keycode[31:24] == 8'h04));
    assign d = ((keycode[15:8] == 8'h07) | (keycode[7:0] == 8'h07)|(keycode[23:16] == 8'h07) | (keycode[31:24] == 8'h07));
    assign w = ((keycode[15:8] == 8'h1A) | (keycode[7:0] == 8'h1A)|(keycode[23:16] == 8'h1A) | (keycode[31:24] == 8'h1A));
    assign s = ((keycode[15:8] == 8'h16) | (keycode[7:0] == 8'h16)|(keycode[23:16] == 8'h16) | (keycode[31:24] == 8'h16));

    mario_image m_i(.*);
    mario_movem m_m(.*);

    always_comb
    begin
        if (mario_x < process + DrawX && DrawX + process < mario_x + 10'd26 && DrawY > mario_y && DrawY < mario_y + 10'd32)
            begin
                mario = 1'b1;
            end
        else
            mario = 1'b0;
    end

endmodule 


module mario_movem (
        input Clk, Reset, frame_clk,
        input w, s, a, d,
        input mario_alive,
        output logic [23:0] mario_counter,
        output logic [9:0] mario_x, mario_y, process, mario_y_motion,
        output logic mario_in_air,
        output logic sl, sr, rr1, rr2, rr3, rl1, rl2, rl3, jr, jl, il, ir, gr, gl, di
);

    parameter [9:0] mario_x_ori = 20;
    parameter [9:0] mario_y_ori = 400;

    parameter [9:0] mario_x_min = 0;
    parameter [9:0] mario_x_max = 639;
    parameter [9:0] mario_y_min = 0;
    parameter [9:0] mario_y_max = 479;
    parameter [9:0] mario_x_step = 2;

    parameter [9:0] mario_x_size = 26;

    logic [9:0] mario_x_motion, level;
    logic [9:0] mario_x_pos_input, mario_x_motion_input, mario_y_pos_input, mario_y_motion_input;
    logic [9:0] process_input;

    logic sl_in, sr_in, rr1_in, rr2_in, rr3_in, rl1_in, rl2_in, rl3_in, jr_in, jl_in, ir_in, il_in, gr_in, gl_in, di_in;

    logic [23:0]  mario_counter_in;
    logic [23:0] counter2, counter2_in;
    logic flag, flag_in;
	logic i;
    always_comb
    begin
        if (mario_y + mario_y_motion >= 10'd384)
            begin
                mario_in_air = 1'b0;
                level = 10'd384;
            end
        else
            begin
                mario_in_air = 1'b1;
                level = 10'd384;
            end
    end

    enum logic [3:0] {STAND_R,
                      STAND_L, 
                      RUN_1_R, 
                      RUN_2_R, 
                      RUN_3_R,
					  RUN_1_L, 
                      RUN_2_L, 
                      RUN_3_L, 
                      JUMP_R,
                      JUMP_L, 
                      IN_AIR_L,
                      IN_AIR_R, 
                      GLIDE_R,
                      GLIDE_L,
                      DIE} STATE, NEXT_STATE;
    
    logic frame_clk_delayed, frame_clk_rising_edge;
    always_ff @ (posedge Clk) 
    begin
        frame_clk_delayed <= frame_clk;
        frame_clk_rising_edge <= (frame_clk == 1'b1) && (frame_clk_delayed == 1'b0);
    end

    always_ff @ (posedge Clk)
    begin
        if (Reset)
            begin
                mario_x <= 10'd80;
                mario_y <= 10'd384;
                mario_x_motion <= 10'd0;
                mario_y_motion <= 10'd0;
                process <= 10'd0;
                STATE <= STAND_R;
                mario_counter <= 24'b0;
                counter2 <= 24'b0;
                flag <= 1'b0;
                sr  <= 1'b1;
                sl  <= 1'b0;
                rr1 <= 1'b0;
                rr2 <= 1'b0; 
                rr3 <= 1'b0; 
                rl1 <= 1'b0; 
                rl2 <= 1'b0; 
                rl3 <= 1'b0; 
                jr  <= 1'b0; 
                jl  <= 1'b0;
                ir  <= 1'b0;
                il  <= 1'b0; 
                gr  <= 1'b0;
                gl  <= 1'b0;
                di  <= 1'b0;
            end
        else
            begin
                mario_x <= mario_x_pos_input;
                mario_y <= mario_y_pos_input;
                mario_x_motion <= mario_x_motion_input;
                mario_y_motion <= mario_y_motion_input;
                process <= process_input;
                STATE <= NEXT_STATE;
                mario_counter <= mario_counter_in;
                counter2 <= counter2_in;
                flag <= flag_in;
                sr  <= sr_in;
                sl  <= sl_in;
                rr1 <= rr1_in;
                rr2 <= rr2_in; 
                rr3 <= rr3_in; 
                rl1 <= rl1_in; 
                rl2 <= rl2_in; 
                rl3 <= rl3_in; 
                jr  <= jr_in; 
                jl  <= jl_in;
                ir  <= ir_in;
                il  <= il_in; 
                gr  <= gr_in;
                gl  <= gl_in;
                di  <= di_in;
            end
    end

    always_comb
    begin
        mario_x_pos_input = mario_x;
        mario_y_pos_input = mario_y;
        mario_x_motion_input = mario_x_motion;
        mario_y_motion_input = mario_y_motion;
        process_input = process;
        NEXT_STATE = STATE;
        flag_in = flag;
        mario_counter_in = mario_counter;
        counter2_in = counter2;
        if (frame_clk_rising_edge)
            begin
                unique case (STATE)
                    default: 
                        begin
                            sr_in  = 1'b0;
                            sl_in  = 1'b0;
                            rr1_in = 1'b0;
                            rr2_in = 1'b0; 
                            rr3_in = 1'b0; 
                            rl1_in = 1'b0; 
                            rl2_in = 1'b0; 
                            rl3_in = 1'b0; 
                            jr_in  = 1'b0; 
                            jl_in  = 1'b0;
                            ir_in  = 1'b0;
                            il_in  = 1'b0; 
                            gr_in  = 1'b0;
                            gl_in  = 1'b0;
                            di_in  = 1'b0;
                        end

                    STAND_R:
                        begin
                            mario_x_motion_input = 10'd0;
                            mario_y_motion_input = 10'd0;
                            mario_counter_in = 24'b0;
                            counter2_in = 24'b0;
                            sr_in  = 1'b1;
                            sl_in  = 1'b0;
                            rr1_in = 1'b0;
                            rr2_in = 1'b0; 
                            rr3_in = 1'b0; 
                            rl1_in = 1'b0; 
                            rl2_in = 1'b0; 
                            rl3_in = 1'b0; 
                            jr_in  = 1'b0; 
                            jl_in  = 1'b0;
                            ir_in  = 1'b0;
                            il_in  = 1'b0; 
                            gr_in  = 1'b0;
                            gl_in  = 1'b0;
                            di_in  = 1'b0;
                            if (mario_alive == 1'b0)
                                begin
                                    NEXT_STATE = DIE;
                                    mario_x_motion_input = 10'd0;
                                    mario_y_motion_input = ~(10'd15) + 1'd1;
                                end
                            else if (w && ~flag)
                                begin
                                    NEXT_STATE = JUMP_R;
                                    flag_in = 1'b1;
                                end
                            else if (a)
                                begin
                                    NEXT_STATE = RUN_1_L;
                                    flag_in = 1'b0;
                                end
                            else if (d)
                                begin
                                    NEXT_STATE = RUN_1_R;
                                    flag_in = 1'b0;
                                end
                            else if (~w)
                                begin
                                    NEXT_STATE = STAND_R;
                                    flag_in = 1'b0;
                                end
                            else
                                begin
                                    NEXT_STATE = STAND_R;
                                    flag_in = flag;
                                end
                        end
                    
                    STAND_L:
                        begin
                            mario_x_motion_input = 10'd0;
                            mario_y_motion_input = 10'd0;
                            mario_counter_in = 24'b0;
                            counter2_in = 24'b0;
                            sr_in  = 1'b0;
                            sl_in  = 1'b1;
                            rr1_in = 1'b0;
                            rr2_in = 1'b0; 
                            rr3_in = 1'b0; 
                            rl1_in = 1'b0; 
                            rl2_in = 1'b0; 
                            rl3_in = 1'b0; 
                            jr_in  = 1'b0; 
                            jl_in  = 1'b0;
                            ir_in  = 1'b0;
                            il_in  = 1'b0; 
                            gr_in  = 1'b0;
                            gl_in  = 1'b0;
                            di_in  = 1'b0;
                            if (mario_alive == 1'b0)
                                begin
                                    NEXT_STATE = DIE;
                                    mario_x_motion_input = 10'd0;
                                    mario_y_motion_input = ~(10'd15) + 1'd1;
                                end
                            else if (w && ~flag)
                                begin
                                    NEXT_STATE = JUMP_L;
                                    flag_in = 1'b1;
                                end
                            else if (a)
                                begin
                                    NEXT_STATE = RUN_1_L;
                                    flag_in = 1'b0;
                                end
                            else if (d)
                                begin
                                    NEXT_STATE = RUN_1_R;
                                    flag_in = 1'b0;
                                end
                            else if (~w)
                                begin
                                    NEXT_STATE = STAND_L;
                                    flag_in = 1'b0;
                                end
                            else
                                begin
                                    NEXT_STATE = STAND_L;
                                    flag_in = flag;
                                end
                        end
                    
                    RUN_1_R:
                        begin
                            mario_x_motion_input = 10'd2;
                            mario_y_motion_input = 10'd0;
                            flag_in = flag;
                            sr_in  = 1'b0;
                            sl_in  = 1'b0;
                            rr1_in = 1'b1;
                            rr2_in = 1'b0; 
                            rr3_in = 1'b0; 
                            rl1_in = 1'b0; 
                            rl2_in = 1'b0; 
                            rl3_in = 1'b0; 
                            jr_in  = 1'b0; 
                            jl_in  = 1'b0;
                            ir_in  = 1'b0;
                            il_in  = 1'b0; 
                            gr_in  = 1'b0;
                            gl_in  = 1'b0;
                            di_in  = 1'b0;
                            if (mario_x + mario_x_size >= mario_x_max)
                                begin
                                    mario_x_motion_input = 10'd0;
                                end
                            if (~w)
                                begin
                                    flag_in = 1'b0;
                                end
                            if (mario_alive == 1'd0)
                                begin
                                    NEXT_STATE = DIE;
                                    mario_x_motion_input = 10'd0;
                                    mario_y_motion_input = ~(9'd15) + 1'd1;
                                end
                            else if (w && ~flag)
                                begin
                                    NEXT_STATE = JUMP_R;
                                    flag_in = 1'b1;
                                end
                            else if (d && mario_counter[3])
                                begin
                                    NEXT_STATE = RUN_2_R;
                                end
                            else if (d && ~mario_counter[3])
                                begin
                                    NEXT_STATE = RUN_1_R;
                                    if (counter2[3] == 1'b1)
                                        begin
                                            mario_counter_in = mario_counter + 24'b1;
                                            counter2_in = counter2 + 24'b1;
                                        end
                                    else 
                                        begin
                                            mario_counter_in = mario_counter;
                                            counter2_in = counter2 + 24'b1;
                                        end
                                end
                            else 
                                begin
                                    NEXT_STATE = STAND_R;
                                end
                        end

                    RUN_2_R:
                        begin
                            mario_x_motion_input = 10'd2;
                            mario_y_motion_input = 10'd0;
                            flag_in = flag;
                            sr_in  = 1'b0;
                            sl_in  = 1'b0;
                            rr1_in = 1'b0;
                            rr2_in = 1'b1; 
                            rr3_in = 1'b0; 
                            rl1_in = 1'b0; 
                            rl2_in = 1'b0; 
                            rl3_in = 1'b0; 
                            jr_in  = 1'b0; 
                            jl_in  = 1'b0;
                            ir_in  = 1'b0;
                            il_in  = 1'b0; 
                            gr_in  = 1'b0;
                            gl_in  = 1'b0;
                            di_in  = 1'b0;
                            if (mario_x + mario_x_size >= mario_x_max)
                                begin
                                    mario_x_motion_input = 10'd0;
                                end
                            if (~w)
                                begin
                                    flag_in = 1'b0;
                                end
                            if (mario_alive == 1'd0)
                                begin
                                    NEXT_STATE = DIE;
                                    mario_x_motion_input = 10'd0;
                                    mario_y_motion_input = ~(10'd15) + 1'd1;
                                end
                            else if (w && ~flag)
                                begin
                                    NEXT_STATE = JUMP_R;
                                    flag_in = 1'b1;
                                end
                            else if (d && mario_counter[3])
                                begin
                                    NEXT_STATE = RUN_3_R;
                                end
                            else if (d && ~mario_counter[3])
                                begin
                                    NEXT_STATE = RUN_2_R;
                                    if (counter2[3] == 1'b1)
                                        begin
                                            mario_counter_in = mario_counter + 24'b1;
                                            counter2_in = counter2 + 24'b1;
                                        end
                                    else 
                                        begin
                                            mario_counter_in = mario_counter;
                                            counter2_in = counter2 + 24'b1;
                                        end
                                end
                            else 
                                begin
                                    NEXT_STATE = STAND_R;
                                end
                        end

                    RUN_3_R:
                        begin
                            mario_x_motion_input = 10'd2;
                            mario_y_motion_input = 10'd0;
                            flag_in = flag;
                            sr_in  = 1'b0;
                            sl_in  = 1'b0;
                            rr1_in = 1'b0;
                            rr2_in = 1'b0; 
                            rr3_in = 1'b1; 
                            rl1_in = 1'b0; 
                            rl2_in = 1'b0; 
                            rl3_in = 1'b0; 
                            jr_in  = 1'b0; 
                            jl_in  = 1'b0;
                            ir_in  = 1'b0;
                            il_in  = 1'b0; 
                            gr_in  = 1'b0;
                            gl_in  = 1'b0;
                            di_in  = 1'b0;
                            if (mario_x + mario_x_size >= mario_x_max)
                                begin
                                    mario_x_motion_input = 10'd0;
                                end
                            if (~w)
                                begin
                                    flag_in = 1'b0;
                                end
                            if (mario_alive == 1'd0)
                                begin
                                    NEXT_STATE = DIE;
                                    mario_x_motion_input = 10'd0;
                                    mario_y_motion_input = ~(10'd15) + 1'd1;
                                end
                            else if (w && ~flag)
                                begin
                                    NEXT_STATE = JUMP_R;
                                    flag_in = 1'b1;
                                end
                            else if (d && mario_counter[3])
                                begin
                                    NEXT_STATE = RUN_1_R;
                                end
                            else if (d && ~mario_counter[3])
                                begin
                                    NEXT_STATE = RUN_3_R;
                                    if (counter2[3] == 1'b1)
                                        begin
                                            mario_counter_in = mario_counter + 24'b1;
                                            counter2_in = counter2 + 24'b1;
                                        end
                                    else 
                                        begin
                                            mario_counter_in = mario_counter;
                                            counter2_in = counter2 + 24'b1;
                                        end
                                end
                            else 
                                begin
                                    NEXT_STATE = STAND_R;
                                end
                        end

                    RUN_1_L:
                        begin
                            mario_x_motion_input = (~10'd2) + 1'b1;
                            mario_y_motion_input = 10'd0;
                            flag_in = flag;
                            sr_in  = 1'b0;
                            sl_in  = 1'b0;
                            rr1_in = 1'b0;
                            rr2_in = 1'b0; 
                            rr3_in = 1'b0; 
                            rl1_in = 1'b1; 
                            rl2_in = 1'b0; 
                            rl3_in = 1'b0; 
                            jr_in  = 1'b0; 
                            jl_in  = 1'b0;
                            ir_in  = 1'b0;
                            il_in  = 1'b0; 
                            gr_in  = 1'b0;
                            gl_in  = 1'b0;
                            di_in  = 1'b0;
                            if (mario_x + mario_x_motion <= 10'd1)
                                begin
                                    mario_x_motion_input = 10'd0;
                                end
                            if (~w)
                                begin
                                    flag_in = 1'b0;
                                end
                            if (mario_alive == 1'd0)
                                begin
                                    NEXT_STATE = DIE;
                                    mario_x_motion_input = 10'd0;
                                    mario_y_motion_input = ~(10'd15) + 1'd1;
                                end
                            else if (w && ~flag)
                                begin
                                    NEXT_STATE = JUMP_L;
                                    flag_in = 1'b1;
                                end
                            else if (a && mario_counter[3])
                                begin
                                    NEXT_STATE = RUN_2_L;
                                end
                            else if (a && ~mario_counter[3])
                                begin
                                    NEXT_STATE = RUN_1_L;
                                    if (counter2[3] == 1'b1)
                                        begin
                                            mario_counter_in = mario_counter + 24'b1;
                                            counter2_in = counter2 + 24'b1;
                                        end
                                    else 
                                        begin
                                            mario_counter_in = mario_counter;
                                            counter2_in = counter2 + 24'b1;
                                        end
                                end
                            else 
                                begin
                                    NEXT_STATE = STAND_L;
                                end
                        end
                    
                    RUN_2_L:
                        begin
                            mario_x_motion_input = (~10'd2) + 1'b1;
                            mario_y_motion_input = 10'd0;
                            flag_in = flag;
                            sr_in  = 1'b0;
                            sl_in  = 1'b0;
                            rr1_in = 1'b0;
                            rr2_in = 1'b0; 
                            rr3_in = 1'b0; 
                            rl1_in = 1'b0; 
                            rl2_in = 1'b1; 
                            rl3_in = 1'b0; 
                            jr_in  = 1'b0; 
                            jl_in  = 1'b0;
                            ir_in  = 1'b0;
                            il_in  = 1'b0; 
                            gr_in  = 1'b0;
                            gl_in  = 1'b0;
                            di_in  = 1'b0;
                            if (mario_x + mario_x_motion <= 10'd1)
                                begin
                                    mario_x_motion_input = 10'd0;
                                end
                            if (~w)
                                begin
                                    flag_in = 1'b0;
                                end
                            if (mario_alive == 1'd0)
                                begin
                                    NEXT_STATE = DIE;
                                    mario_x_motion_input = 10'd0;
                                    mario_y_motion_input = ~(10'd15) + 1'd1;
                                end
                            else if (w && ~flag)
                                begin
                                    NEXT_STATE = JUMP_L;
                                    flag_in = 1'b1;
                                end
                            else if (a && mario_counter[3])
                                begin
                                    NEXT_STATE = RUN_3_L;
                                end
                            else if (a && ~mario_counter[3])
                                begin
                                    NEXT_STATE = RUN_2_L;
                                    if (counter2[3] == 1'b1)
                                        begin
                                            mario_counter_in = mario_counter + 24'b1;
                                            counter2_in = counter2 + 24'b1;
                                        end
                                    else 
                                        begin
                                            mario_counter_in = mario_counter;
                                            counter2_in = counter2 + 24'b1;
                                        end
                                end
                            else 
                                begin
                                    NEXT_STATE = STAND_L;
                                end
                        end
                    
                    RUN_3_L:
                        begin
                            mario_x_motion_input = (~10'd2) + 1'b1;
                            mario_y_motion_input = 10'd0;
                            flag_in = flag;
                            sr_in  = 1'b0;
                            sl_in  = 1'b0;
                            rr1_in = 1'b0;
                            rr2_in = 1'b0; 
                            rr3_in = 1'b0; 
                            rl1_in = 1'b0; 
                            rl2_in = 1'b0; 
                            rl3_in = 1'b1; 
                            jr_in  = 1'b0; 
                            jl_in  = 1'b0;
                            ir_in  = 1'b0;
                            il_in  = 1'b0; 
                            gr_in  = 1'b0;
                            gl_in  = 1'b0;
                            di_in  = 1'b0;
                            if (mario_x + mario_x_motion <= 10'd1)
                                begin
                                    mario_x_motion_input = 10'd0;
                                end
                            if (~w)
                                begin
                                    flag_in = 1'b0;
                                end
                            if (mario_alive == 1'd0)
                                begin
                                    NEXT_STATE = DIE;
                                    mario_x_motion_input = 10'd0;
                                    mario_y_motion_input = ~(10'd15) + 1'd1;
                                end
                            else if (w && ~flag)
                                begin
                                    NEXT_STATE = JUMP_L;
                                    flag_in = 1'b1;
                                end
                            else if (a && mario_counter[3])
                                begin
                                    NEXT_STATE = RUN_1_L;
                                end
                            else if (a && ~mario_counter[3])
                                begin
                                    NEXT_STATE = RUN_3_L;
                                    if (counter2[3] == 1'b1)
                                        begin
                                            mario_counter_in = mario_counter + 24'b1;
                                            counter2_in = counter2 + 24'b1;
                                        end
                                    else 
                                        begin
                                            mario_counter_in = mario_counter;
                                            counter2_in = counter2 + 24'b1;
                                        end
                                end
                            else 
                                begin
                                    NEXT_STATE = STAND_L;
                                end
                        end
                    
                    JUMP_R:
                        begin
                            sr_in  = 1'b0;
                            sl_in  = 1'b0;
                            rr1_in = 1'b0;
                            rr2_in = 1'b0; 
                            rr3_in = 1'b0; 
                            rl1_in = 1'b0; 
                            rl2_in = 1'b0; 
                            rl3_in = 1'b0; 
                            jr_in  = 1'b1; 
                            jl_in  = 1'b0;
                            ir_in  = 1'b0;
                            il_in  = 1'b0; 
                            gr_in  = 1'b0;
                            gl_in  = 1'b0;
                            di_in  = 1'b0;
                            mario_x_motion_input = mario_x_motion;
                            mario_y_motion_input = (~10'd15) + 1'd1;
                            flag_in = 1'b1;
                            NEXT_STATE = IN_AIR_R;
                        end
                    
                    JUMP_L:
                        begin
                            sr_in  = 1'b0;
                            sl_in  = 1'b0;
                            rr1_in = 1'b0;
                            rr2_in = 1'b0; 
                            rr3_in = 1'b0; 
                            rl1_in = 1'b0; 
                            rl2_in = 1'b0; 
                            rl3_in = 1'b0; 
                            jr_in  = 1'b0; 
                            jl_in  = 1'b1;
                            ir_in  = 1'b0;
                            il_in  = 1'b0; 
                            gr_in  = 1'b0;
                            gl_in  = 1'b0;
                            di_in  = 1'b0;
                            mario_x_motion_input = mario_x_motion;
                            mario_y_motion_input = (~10'd15) + 1'd1;
                            flag_in = 1'b1;
                            NEXT_STATE = IN_AIR_L;
                        end
                    
                    IN_AIR_R:
                        begin
                            sr_in  = 1'b0;
                            sl_in  = 1'b0;
                            rr1_in = 1'b0;
                            rr2_in = 1'b0; 
                            rr3_in = 1'b0; 
                            rl1_in = 1'b0; 
                            rl2_in = 1'b0; 
                            rl3_in = 1'b0; 
                            jr_in  = 1'b0; 
                            jl_in  = 1'b0;
                            ir_in  = 1'b1;
                            il_in  = 1'b0; 
                            gr_in  = 1'b0;
                            gl_in  = 1'b0;
                            di_in  = 1'b0;
                            if (a && ~d && mario_x_motion_input == 10'd0)
                                begin
                                    mario_x_motion_input = (~10'd2) + 1'b1;
        
                                    if (mario_x + mario_x_motion_input <= 10'd1)
                                        begin
                                            mario_x_motion_input = 10'd0;
                                        end
                                end
                            else if (~a && d && mario_x_motion_input == 10'd0)
                                begin
                                    mario_x_motion_input = 10'd2;
                                    if (mario_x + mario_x_motion_input >= 10'd439)
                                        begin
                                            mario_x_motion_input = 10'd0;
                                        end
                                end
                            else
                                begin
                                    mario_x_motion_input = mario_x_motion;
                                end

                            flag_in = 1'b1;
                            if (mario_alive == 1'b0)
                                begin
                                    NEXT_STATE = DIE;
                                    mario_x_motion_input = 10'd0;
                                    mario_y_motion_input = ~(10'd15) + 1'd1;
                                end
                            else
                                begin
                                    if (mario_in_air)
                                        begin
                                            NEXT_STATE = IN_AIR_R;
                                            mario_y_motion_input = mario_y_motion + 1'd1;
                                            if (mario_y + mario_y_motion < 10'd5)
                                                begin
                                                    mario_y_motion_input = (~mario_y_motion) + 10'd1;
                                                end
                                        end
                                    else
                                        begin
                                            if (a == 1'b1)
                                                begin
                                                    NEXT_STATE = GLIDE_L;
                                                end
                                            else 
                                                begin
                                                    NEXT_STATE = GLIDE_R;
                                                end
                                            mario_y_motion_input = 10'd0;
                                            if (w)
                                                begin
                                                    flag_in = 1'b1;
                                                end
                                            else
                                                begin
                                                    flag_in = 1'b0;
                                                end
                                        end
                                end
                        end

                    IN_AIR_L:
                        begin
                            sr_in  = 1'b0;
                            sl_in  = 1'b0;
                            rr1_in = 1'b0;
                            rr2_in = 1'b0; 
                            rr3_in = 1'b0; 
                            rl1_in = 1'b0; 
                            rl2_in = 1'b0; 
                            rl3_in = 1'b0; 
                            jr_in  = 1'b0; 
                            jl_in  = 1'b0;
                            ir_in  = 1'b0;
                            il_in  = 1'b1; 
                            gr_in  = 1'b0;
                            gl_in  = 1'b0;
                            di_in  = 1'b0;
                            if (a && ~d && mario_x_motion_input == 10'd0)
                                begin
                                    mario_x_motion_input = (~10'd2) + 1'b1;
        
                                    if (mario_x + mario_x_motion_input <= 10'd1)
                                        begin
                                            mario_x_motion_input = 10'd0;
                                        end
                                end
                            else if (~a && d && mario_x_motion_input == 10'd0)
                                begin
                                    mario_x_motion_input = 10'd2;
                                    if (mario_x + mario_x_motion_input >= 10'd439)
                                        begin
                                            mario_x_motion_input = 10'd0;
                                        end
                                end
                            else
                                begin
                                    mario_x_motion_input = mario_x_motion;
                                end

                            flag_in = 1'b1;
                            if (mario_alive == 1'b0)
                                begin
                                    NEXT_STATE = DIE;
                                    mario_x_motion_input = 10'd0;
                                    mario_y_motion_input = ~(10'd15) + 1'd1;
                                end
                            else
                                begin
                                    if (mario_in_air)
                                        begin
                                            NEXT_STATE = IN_AIR_L;
                                            mario_y_motion_input = mario_y_motion + 1'd1;
                                            if (mario_y + mario_y_motion < 10'd5)
                                                begin
                                                    mario_y_motion_input = (~mario_y_motion) + 10'd1;
                                                end
                                        end
                                    else
                                        begin
                                            if (a == 1'b1)
                                                begin
                                                    NEXT_STATE = GLIDE_L;
                                                end
                                            else 
                                                begin
                                                    NEXT_STATE = GLIDE_R;
                                                end
                                            mario_y_motion_input = 10'd0;
                                            if (w)
                                                begin
                                                    flag_in = 1'b1;
                                                end
                                            else
                                                begin
                                                    flag_in = 1'b0;
                                                end
                                        end
                                end
                        end
                    
                    GLIDE_R:
                        begin
                            mario_x_motion_input = mario_x_motion;
                            sr_in  = 1'b0;
                            sl_in  = 1'b0;
                            rr1_in = 1'b0;
                            rr2_in = 1'b0; 
                            rr3_in = 1'b0; 
                            rl1_in = 1'b0; 
                            rl2_in = 1'b0; 
                            rl3_in = 1'b0; 
                            jr_in  = 1'b0; 
                            jl_in  = 1'b0;
                            ir_in  = 1'b0;
                            il_in  = 1'b0; 
                            gr_in  = 1'b1;
                            gl_in  = 1'b0;
                            di_in  = 1'b0;
                            if (mario_alive == 1'd0)
                                begin
                                    NEXT_STATE = DIE;
                                    mario_x_motion_input = 10'd0;
                                    mario_y_motion_input = ~(10'd15) + 1'd1;
                                end
                            else if (mario_x + mario_x_size >= mario_x_max)
                                begin
                                    mario_x_motion_input = 10'd0;
                                end
                            else if (mario_x <= process + 10'd0)
                                begin
                                    mario_x_motion_input = 10'd0;
                                end
                            else
                                begin
                                    if (mario_x_motion == 10'd0)
                                        begin
                                            NEXT_STATE = STAND_R;
                                        end
                                    else if (mario_x_motion == 10'd1)
                                        begin
                                            NEXT_STATE = RUN_1_R;
                                        end
                                    else if (mario_x_motion == 10'd2)
                                        begin
                                            NEXT_STATE = RUN_2_R;
                                        end
                                    else if (mario_x_motion == 10'd3)
                                        begin
                                            NEXT_STATE = RUN_3_R;
                                        end
                                    else if (mario_x_motion == (~10'd1) + 1'b1)
                                        begin
                                            NEXT_STATE = RUN_1_L;
                                        end
                                    else if (mario_x_motion == (~10'd2) + 1'b1)
                                        begin
                                            NEXT_STATE = RUN_2_L;
                                        end
                                    else if (mario_x_motion == (~10'd3) + 1'b1)
                                        begin
                                            NEXT_STATE = RUN_3_L;
                                        end
                                    else
                                        NEXT_STATE = STAND_R;
                                end
                        end

                    GLIDE_L:
                        begin
                            mario_x_motion_input = mario_x_motion;
                            sr_in  = 1'b0;
                            sl_in  = 1'b0;
                            rr1_in = 1'b0;
                            rr2_in = 1'b0; 
                            rr3_in = 1'b0; 
                            rl1_in = 1'b0; 
                            rl2_in = 1'b0; 
                            rl3_in = 1'b0; 
                            jr_in  = 1'b0; 
                            jl_in  = 1'b0;
                            ir_in  = 1'b0;
                            il_in  = 1'b0; 
                            gr_in  = 1'b0;
                            gl_in  = 1'b1;
                            di_in  = 1'b0;
                            if (mario_alive == 1'd0)
                                begin
                                    NEXT_STATE = DIE;
                                    mario_x_motion_input = 10'd0;
                                    mario_y_motion_input = ~(10'd15) + 1'd1;
                                end
                            else if (mario_x + mario_x_size >= mario_x_max)
                                begin
                                    mario_x_motion_input = 10'd0;
                                end
                            else if (mario_x <= process + 10'd0)
                                begin
                                    mario_x_motion_input = 10'd0;
                                end
                            else
                                begin
                                    if (mario_x_motion == 10'd0)
                                        begin
                                            NEXT_STATE = STAND_L;
                                        end
                                    else if (mario_x_motion == 10'd1)
                                        begin
                                            NEXT_STATE = RUN_1_R;
                                        end
                                    else if (mario_x_motion == 10'd2)
                                        begin
                                            NEXT_STATE = RUN_2_R;
                                        end
                                    else if (mario_x_motion == 10'd3)
                                        begin
                                            NEXT_STATE = RUN_3_R;
                                        end
                                    else if (mario_x_motion == (~10'd1) + 1'b1)
                                        begin
                                            NEXT_STATE = RUN_1_L;
                                        end
                                    else if (mario_x_motion == (~10'd2) + 1'b1)
                                        begin
                                            NEXT_STATE = RUN_2_L;
                                        end
                                    else if (mario_x_motion == (~10'd3) + 1'b1)
                                        begin
                                            NEXT_STATE = RUN_3_L;
                                        end
                                    else
                                        NEXT_STATE = STAND_L;
                                end
                        end
                    
                    DIE:
                        begin
                            sr_in  = 1'b0;
                            sl_in  = 1'b0;
                            rr1_in = 1'b0;
                            rr2_in = 1'b0; 
                            rr3_in = 1'b0; 
                            rl1_in = 1'b0; 
                            rl2_in = 1'b0; 
                            rl3_in = 1'b0; 
                            jr_in  = 1'b0; 
                            jl_in  = 1'b0;
                            ir_in  = 1'b0;
                            il_in  = 1'b0; 
                            gr_in  = 1'b0;
                            gl_in  = 1'b0;
                            di_in  = 1'b1;
                            NEXT_STATE = DIE;
                            mario_y_motion_input = mario_y_motion + 1'd1;
                        end
                endcase
                
                mario_x_pos_input = mario_x + mario_x_motion;
                if (mario_x_pos_input >= mario_x_max)
                    begin
                        mario_x_pos_input = mario_x_max;
                    end
                if (mario_in_air || (STATE == DIE))
                    begin
                        mario_y_pos_input = mario_y + mario_y_motion;
                        if ((STATE == DIE) && (mario_y + mario_y_motion >= mario_y_max))
                            begin
                                mario_y_pos_input = mario_y_max;
                            end
                    end
                else
                    begin
                        mario_y_pos_input = level;
                    end
            end
        else
            begin
                sr_in  = sr;
                sl_in  = sl;
                rr1_in = rr1;
                rr2_in = rr2; 
                rr3_in = rr3; 
                rl1_in = rl1; 
                rl2_in = rl2; 
                rl3_in = rl3; 
                jr_in  = jr; 
                jl_in  = jl;
                ir_in  = ir;
                il_in  = il; 
                gr_in  = gr;
                gl_in  = gl;
                di_in  = di;
            end
    end
endmodule
                
module mario_image (
        input Clk, Reset, frame_clk,
        input [9:0] mario_x,
        input sl, sr, rr1, rr2, rr3, rl1, rl2, rl3, jr, jl, ir, gr, gl, di,il,
        input [23:0] mario_sl, mario_sr, mario_rl1, mario_rl2, mario_rl3, mario_rr1, mario_rr2, mario_rr3, mario_jr, mario_jl, mario_die,
        output [23:0] mario_pic_out
);
    always_ff @ (posedge Clk)
        begin
            if (sl == 1'b1)
                begin
                    mario_pic_out = mario_sl;
                end
            else if (sr == 1'b1)
                begin
                    mario_pic_out = mario_sr;
                end
            else if (rr1 == 1'b1)
                begin
                    mario_pic_out = mario_rr1;
                end
            else if (rr2 == 1'b1)
                begin
                    mario_pic_out = mario_rr2;
                end
            else if (rr3 == 1'b1)
                begin
                    mario_pic_out = mario_rr3;
                end
            else if (rl1 == 1'b1)
                begin
                    mario_pic_out = mario_rl1;
                end
            else if (rl2 == 1'b1)
                begin
                    mario_pic_out = mario_rl2;
                end
            else if (rl3 == 1'b1)
                begin
                    mario_pic_out = mario_rl3;
                end
            else if (jr == 1'b1)
                begin
                    mario_pic_out = mario_jr;
                end
            else if (jl == 1'b1)
                begin
                    mario_pic_out = mario_jl;
                end
            else if (ir == 1'b1)
                begin
                    mario_pic_out = mario_jr;
                end
            else if (il == 1'b1)
                begin
                    mario_pic_out = mario_jl;
                end
            else if (gr == 1'b1)
                begin
                    mario_pic_out = mario_jr;
                end
            else if (gl == 1'b1)
                begin
                    mario_pic_out = mario_jl;
                end
            else if (di == 1'b1)
                begin
                    mario_pic_out = mario_die;
                end
            else
                begin
                    mario_pic_out = mario_sr;
                end
            
        end
    
endmodule