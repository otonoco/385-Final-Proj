    Mac OS X            	   2   �                                           ATTR         �   L                  �     com.apple.lastuseddate#PS       �   <  com.apple.quarantine ձ_    j�^    q/0083;5fb1d05b;Safari;CBE46DCC-8259-4AAD-823C-D8AAEC365727 