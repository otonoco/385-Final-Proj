    Mac OS X            	   2  y     �                                      ATTR      �  @  k                 @     com.apple.lastuseddate#PS      P   H  com.apple.macl     �   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms   o   <  com.apple.quarantine �u�_    �Y�8     �x9(8�CѸ�C�5-�                                                       bplist00�3A¬��Y�"
                            bplist00�_shttps://wiki.illinois.edu/wiki/download/attachments/728156926/font_rom.sv?version=1&modificationDate=1596810123000&
                            �q/0083;5fa9b3c0;Safari;3E43F65C-F436-4B97-BB6C-CA3963555436 